module fifo(clk,rst,wdata,rdata,wr_en,rd_en,full,empty);
input clk,rst,wr_en,rd_en;
output full,empty;
  input [7:0] wdata;
  output reg [7:0] rdata;

  reg [5:0] wr_ptr;
  reg [5:0] rd_ptr;

reg [7:0]mem[31:0];

integer i;
//writing data into fifo
always @(posedge clk,posedge rst)
    if (rst) begin

        for(i=0;i<32;i=i+1)
            mem[i]<=8'b0;
         //  wr_ptr<=1'b0;
            end

    else if (wr_en & ~full)
      //mem[{wr_ptr[4],wr_ptr[3],wr_ptr[2],wr_ptr[1],wr_ptr[0]}]<=wdata;
      mem [wr_ptr]<=wdata;


 //reading from fifo
always @(posedge clk,posedge rst)
    if(rst) begin

           //  rd_ptr=1'b0;
             rdata<=8'b0;
         end

    else if (rd_en & ~empty)
        //rdata<=mem[{rd_ptr[4],rd_ptr[3],rd_ptr[2],rd_ptr[1],rd_ptr[0]}];
      rdata<=mem[rd_ptr];

//generating write pointer    
always @(posedge clk,posedge rst)
        if(rst)
            wr_ptr<=6'b0;
        else if(wr_en & ~full)
            wr_ptr<=wr_ptr+1;


always @(posedge clk,posedge rst)
        if(rst)
            rd_ptr<=6'b0;
        else if(rd_en & ~empty)
            rd_ptr<=rd_ptr+1;

assign empty =(rd_ptr==wr_ptr);

assign full=((wr_ptr[4:0]==rd_ptr[4:0])&&(wr_ptr[5]!=rd_ptr[5]));

endmodule
